// 数据存储器
module dm(
    Ad,WrData,DMWr, Clk,
    DM
);
input [31:2] Ad;
input [31:0] WrData;
input DMWr, Clk;
output DM[31:0];

// TODO

endmodule // dm