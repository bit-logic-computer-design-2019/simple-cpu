// 指令存储器，读入一个地址，输出那个地址所存储的数据
module im(
    PC,
    IM
);
input PC[32:2];
output IM[32:0];

// 利用某种方式读取


endmodule //i