module mips(
    
);

endmodule // mips  