module alu(
    A, B,ALUctrl,
    ALU, beq, carrier
);

input [31:0] A;
input [31:0] B;
input ALUctrl[2:0];
output ALU[31:0];
output beq;
output carrier;

// TODO

endmodule // alu  